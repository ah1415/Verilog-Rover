
module atan (
	areset,
	clk,
	q,
	x,
	y);	

	input		areset;
	input		clk;
	output	[8:0]	q;
	input	[11:0]	x;
	input	[11:0]	y;
endmodule
